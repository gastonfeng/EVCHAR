** circuit file for profile: 11 

** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT PROFILES

*Libraries: 
* Local Libraries :
.LIB "D:\my_lib\orcad.lib" 
* From [PSPICE NETLIST] section of pspice91.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500u 0 
.PROBE 
.INC "trans-SCHEMATIC1.net" 

.INC "trans-SCHEMATIC1.als"


.END
